module ldpc_enc(

    );

  
endmodule
