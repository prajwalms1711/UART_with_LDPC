module ldpc_dec(
  );

endmodule
