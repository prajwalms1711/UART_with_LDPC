module ldpc_dec_tb();
endmodule
