module ldpc_enc_tb();
endmodule
